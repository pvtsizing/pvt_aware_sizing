two_stage_amp test

* Two stage OPAMP
.include "../spice_models/gf180/ngspice/design.ngspice"
.lib "../spice_models/gf180/ngspice/sm141064.ngspice" typical

.param wp1=100.0u  lp1=300n mp1=1
.param wn1=8.05u  ln1=300n mn1=1
.param wn3=34.73u ln3=300n mn3=1
.param wp3=7.24u  lp3=300n mp3=1
.param wn4=6.12u  ln4=300n mn4=1
.param wn5=27.11u ln5=300n mn5=1
.param cc=2.95p
.param ibias=30u
.param cload=10p
.param vddh=3.3
.param vcm=0.5*vddh
 


xp1 net4 net4 VDD VDD   pmos_3p3 w=wp1 l=lp1 m=mp1
xp2 net5 net4 VDD VDD   pmos_3p3 w=wp1 l=lp1 m=mp1
xn1 net4 net2 net3 net3 nmos_3p3 w=wn1 l=ln1 m=mn1
xn2 net5 net1 net3 net3 nmos_3p3 w=wn1 l=ln1 m=mn1
xn3 net3 net7 VSS VSS   nmos_3p3 w=wn3 l=ln3 m=mn3
xn4 net7 net7 VSS VSS   nmos_3p3 w=wn4 l=ln4 m=mn4
xp3 net6 net5 VDD VDD   pmos_3p3 w=wp3 l=lp3 m=mp3
xn5 net6 net7 VSS VSS   nmos_3p3 w=wn5 l=ln5 m=mn5
cc net5 net6 {cc}
ibias VDD net7 ibias

vin in 0 dc=0 ac=1.0
ein1 net1 cm in 0 0.5
ein2 net2 cm in 0 -0.5
vcm cm 0 dc=vcm

vdd VDD 0 dc=vddh
vss 0 VSS dc=0
CL net6 0 {cload}


.control
set temp=27
ac dec 10 1 10G
run
set units=degrees
set wr_vecnames
option numdgt=7
wrdata ac.csv v(net6)
op
wrdata dc.csv i(vdd)
dc vin -0.001 0.001 1e-5
wrdata dc_sweep.csv v(net6)
.endc

.end